module fibonocci ( clk, y, reg [3:0] );
  input clk;
  output reg [3:0] y;
               


endmodule
               